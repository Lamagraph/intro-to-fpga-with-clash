../../../src/08-fpga/huffman_top.sv